* resistencias en paralelo
vdd 0 1 vdc=12 type=vdc
vdd1 1 2 vdc=0 type=vdc
vdd2 1 3 vdc=0 type=vdc
vdd3 1 4 vdc=0 type=vdc
r1 2 0 10k
r2 3 0 2k
r3 4 0 1k
.op
.end
